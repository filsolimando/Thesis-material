BZh91AY&SY��� J߀py������?���`�x�4�I��   I�&OB2h     ���#!�4a0F�4b�20 ��!�	�4ѣ4ɑ� �S�AL��h     4 ��!�	�4ѣ4ɑ� �RB@M
`�ԧ�?DOS��82����$�$��~O�JR�����"&ޱ7}�|�d�o���������� �XE$��%ސD��8��|$T��� �Urkݜ@*H�nT6���,�l�-"�{+�L0��kP0�be��.�o�����o�|~^����a�4밌�"6@@����p>�a�KVi3���ّ|_(�FUj�+��L�0z�����ڤ�=[��^�qY[��j8l*WP�TU)�ṽ��ś>����}4u*�_��o[��" ��.�!&��{Fm͊R�4���v�����s�l�t�vGW���ﳊ;"�R��vY�|$eSt���+�S������k����H(�U�Z��j�e\��e�L�k�&>�T�VO#��4o��QT��SU�ӺXq㬹�����&%3g/��nZ����u���v!�+1)S~ۘ�q��Z+��c���6��Y��7�:�@���$a�/[BH4�6�na����LF�!+�i���I�EU*-[M��c:Ýb�3F�M��N3V�3��6巭h��6L�5n�
ZQ��=��$�>�(�.ꪪ��� I'T:�!��#��ؗ���м,R`qw+3yf^KR��j�[�T\�,] �a�6�n��6�fff�b�W�ZؒOʖ�L���*E�{a��
*�iH�Z-R����M8~m�sɷ���� �J�iW�e�Z	����A����B�M�%#d�7�����f��j�n���w����{��}n�XYy�������>6�3��q�㮖|ɳ�+G{(p*��E�3�Gj6���Z�5�m3��;�Z���'�G��i����a�Ls��cRyI�}�i=O�fX��chiαp��'n�0�A���t�b�H���B��a��$��xe���Ny�������#NM�Z����~�V��ƌʌ��Z�rB�T�Eѻ�|���˄X��ǩ9#���E������s��H�k��9��R6�"e��h�d�bz��s���r��v�󲮞9�h�󯤏�NW����4N�W��OgE�'=���G�ɈsL9��?�3m?S>�]l���m�������"u���jEзc��~}�5VN�M�4Lv��G�S���H(���&��Y�mV|���F��2靘��2�80�ڒ�(e�-ͥ�7��$&�*�a��I��2�k�jZ��]Q�г.V�I���V�����0]��Aj���\���;믫��׫��9d��/�Q�y]"�ͽ#��zH~�\}F���w���
�t�^�8�g_G����av�{8aF��F�a�H��UH�t�y�ٗ�~}d��G)3��ng
�Q�E:I��=�m30F��:l��*��>߿d��7q̛rC�T+�94\jF��X�j+H^���ox,�)R�֪Fi��"k�dr�>RN��!vfp����`�zva������*D���N�H��"��Y��Y�EId��������z�"���i�VtҪwK����,�B�<��E��9]����"�(H�wk 