BZh91AY&SYv� 	W_��y���������� @ `{����dZ
 ֐[Z}����Z5#ҁ�4 4�F@   q�&�#F	���h�#@0�OB�� h�      	4�� �P     �A*����j��d4�2M �M4$�B	��M4��&ɦ���A�#&и�1H� B�@�D�C�DD�'�nB�!�G�?���?�Rq���+�_6����X�AFF?�	t�@&[L,�er�
���,!x��H$���/��UZZ��KUUQi%B�0����}W��z��c� =�� �-(G��X���GZg�*9�����'
�ֱ�3]�K"q�)�Q���u��%�P2s�-\h��r%N�D,�	f&�9�ï�U�ob��B�
 ���#r�H0��{uO�V��2�;�d�WX�� �y���<���j�&f��!�5�p*�i��p=��id-�P��ц����vt�%��a�	�9 N�JY�Cp�֝�����!�h�HUT�h!XM��($8MQ&4q,�ѣ��0l�فĶ�ǚ�z�ε���us�LB�_�m��Xd�8�
y6�I*����Hk� Z&�D����6�\�c���y|��i�o��|�O��#��4�Z��ڟey:��$�HH�#/>��C���3�HxI�N�O-��	����k��F��\�I��w���`q�r;L��	��5��&�Qro�c�ck�?��Y�����	4�������vfq��S�K�vĕ�g"TU3H��H��{樔�і6��N�Go��&`kl��-�I����7��%��jN�NJ�R�Øwu�����H�C��[��K)�;s�%w�%h�}a��O6���{a�ɢ�*�g%l)��!s|����;6Y�j�_;�\bҦ.�Nwil�H����'�ݙ=z��$����2�����zo��K�nH�CT���F/���yּ]x	Z�v^�SIۮ��ӓ��c/\�.��;�iۯ�ރ���i4贜��n�����矯�ws�P��N)f:�{K��m�5�38;�c�J���ggSm�r�=��>�{��~�����X"���B��������$�Ib�zWI��Ck�"a3��U;2.1Å�q�emCIcC���ɁΝ'6��m�ner����&��okn.c�k�o[��n�D*f�m\�m�Z嵷+n6���X.Z�?�l!�+R�p���mjr�k>�l�����\5
]�T�T�"i6��U�R"Z7OJ�`222@X� ��f6��߇��\�竫�Ǉ��C[�D��B{�~X�	�v����a�%���̟:}Iꎀ�N�|���$���Ϛ'F���B����M4MH��,jE�:�)�~��fb�$��V�ȝ�$��O�1>�T��BP���J �ԵA,-d+W�s�"w����|?K�,|�?wl�x���b�dP�A��@������i�}\���ʟ)�g܀��@�W�V����$ڝ�db]E��:@�7�|�=�@yE�ʟX�O���JW�x��<�,-�a�g�|[��ҟ���F��&C���������TH�!aA��N��!���)B�'�P�$��"sK�--�VKg�L�P�����z����˿���Ӄv�0P�l)�֡=�,��.Y 6	�Pߺ�8�Zbi��,y��&)�7������8
e�R$�$�!����ډ��d�#�A�E�؜\�pJQ�X7���݂����M�.�N~�8���<�o�~'�Z�N���
]B���lޮ���S^FII{w"}���.�=������ƭ9���y��"�:o��	���L���2�4"]3#��biy�`q!��Y8���[�C�F�݉����؜��չw��2;a%�� �B���1���-�+��8��рj�d��(R��-<�qLB�̱"���D�JD�IJ�~[�J0+������C� ������$/�ҖP����D%&;�A��B�`*0T��4�n � ��覄9�Ɠ�אE��a,J��ڡBy�d�'�]A�Zhĉf��ݡ�cK�U���Pф\�C�C�b�"@"@��s��������>�8籷ω��	�ԛD�Rh)��:3:6P�0�.�BJ�L�OB\?O��I�=���z�ف9"XD���hN]'��	=Ju(U
�Z�=#�&I��&*`�x�
em�hbM���މ�JD���L��	�)Jz��b �D�5�J���i�$�L���5"m��@�Bʀ�J)(��"�Nct��AB���q�p[��Z~��'r[�6!�C5;S�-ޡ��׫�1��8��C,�jP�(d��*��f�%�(�M6�����)��K@`��W�����,X��"6�22i�1�,�P�@K �M�t6S�O[o@D�=	�(@|�6��S�n�e���J ��}�xbŊ�X���(��pw1��ԟA����sD��0���b"Y{��y&C�C����{U�y�<|i�r�{��>F��.�BY�(D�R)C�3����7!_������"�(H;
E 