BZh91AY&SYi��< �_�py����������`	_o5фA]��@P�I�14�i�4���4 �$�i�&�I��L��`bm#�=@=!�M21M0�&�F	���#C@$"h�OSS��4z��2   4�#��i�`��244RDD�ɩ��hFFI��I��1dm�"��JI@�Aɤ���U<��$�I�$:���Tr��<�_�b�	�GF�W��c',��r�1��b��Q�F���Y��m�ߠl#m�;_��lt&����8�A�e���j�d����j"_����0H��H���d=l�Hm�c�9�k�&��K�¶%��(�&*
�C�*v(/����>"~�S(=��a�W��auX���rHˍ6�nu�e^�gn�,�q���wK��8���s{��@3`!��JfOw�
M�V��z�%�U"��K�������Z�a3N��{^��mxV�@�F�*��~lH���V��mى\���9���8ךS9�p}jOφ{���=�ݻ��P��)*��Lex�	g�3�>B�DOS�Jw{��K
K�.`4�Y�-ˬ�㎞2��i`��~f0���b�ͬ-���	�f���k�����)���$����{�H/ q�%c���cB�00̎��`�@�w����m+���w�N���ܽ*H�2hm#�\�޸/qE�ڍ�	��V����!���M�Mol<�J�Thʥ��K���6g5�o�+��������n��<�t�z޴���JU*]5T�m��m��H�=œź�"�+l�ZZ��Xv�[X�L&�E(��I��L�����n�l�F��f*�ނ!l���e�q�Tr��X��#�ʧ�ө2K"��/C!�(�<�2jZ��#*��I��T��)��n�y tS�c�>y�m����S���;�,����)mcV�l�O*F�2�x@��Wew��#):�g����ctd�Iar�m<N��>~�с��+	v�:���k٫���/[9Uz�T���$v�u�5������߾:�|�:�b*G�)(�G��CF��X��K��y�8~ZD�îE�6?��MD��=�c�����|�'���䯕�������K��o�F'��R�L5a��ZӜ��e�Z9��ˌM�4!�b�H�T��eBд=�պF���[�y٫��Rsu7��9>W螬�_vl��NW'6B�W��F2��5�h� ��� 4��B����Ga�.�Չ��66�����"�W���Fhb��	�E>#N=қ���s-o���H��T�MLƄ��<��~�����Ӟ~�P��e�MՄ���nL��7��F��u{Z��Ʒc/�KD�����D{:�<�苰e<m?���v^V�:���E]w%���lss�q�ٱ��ܝ�=�s�I*���-B�[�rd��]�1W��4���w�r8,L�8�Y���Q�v*�P��jF���M)K6�dU!b[��n���iXeücA6�I�FM�FQ�8�F�z��-sV.�"REE�ǝ��X�E"��&���QyER,P���u�A��q�B��Qc#E��A���)
�C4=̒Y�J,�vk�<Ô���Ί���lɰɲ��d��,��O��X��`���6����;\�lU"�$`���Uq�wwEP�G������K�!��S��5_�T�s>G��Q��#�1�u���v2�թ��򅡱���~�[#&,�mmB�"�h�Y��I�0R���v/!ukG��u/�M%l푤*Y՞߶a"g��bM&�/�1�N�><��fV��ۺ��ѪB֗InH��o�31cc��4Ø��!t�v�R�Dᡵ�04lt�ƸT�MEګ����7i݌�RE&�a��n��$�q|`ޑ�2�o1gO���`*�*�N\�Ux�洏�`s�N�|���":�|�OYQP�=��є���ܑN$a1� 