BZh91AY&SY�/�' M_��y������?���@   `�W�����U��0*@6�J�%1O&���MOD4 �z�� d*���@      i���i��4�0LL�������4 h     ���h����h�F@� � �A$ɲ*6��Sj4i�� ��4�dԂ����?�!B!�*�!1�;����B��b�8[�<���D{�-�A�E� �������u   �.�LP�`VZ���%����LVT�6�D2��J�&,�QUuSmj#��e
�,d�Y;�J�f�n����8F^ō�{�j8�#u���lcbA���9��^�E�Y'����~%�h�»�oY%�V�=�(+�+[��*�^�g�P+&I�������ya�N<n]q/�h'`xA�$٨�.	f��'��v�BM곅ܲ���i��U�7�YU�����D9�=G�J
��II�|(��3�1�a"%&H8p� ��H��80KfIk�c��'GF����a��ܫ�B�5��MtM�,�\+�b"V�J,EЪ�+�((FR��F١����GV8
���҆J������ݻ@�;��rb�l��&nX"%A����2�sV��J�t��)5��,��8��Ǝ%�i�[�`�[��#��7qe��e6M����Zԃ����69�V�N��#=��7$���hR��3*������,%�R�f^*�+JT=!*����*u7=g7���t9���I����e_+��/_��z�p��A ��-�      � �Q�O=A�>����68���b�$�u�Q[`��%����]�¦y]�Wu$����.�$�(Ks\Ҍm6�@��44H]�R�D@}��bT h.q���!"�-p��$�`��K�]�f�������F��W#�?=�e`E��ÈF�&On�:K(V*U\*��$q/!
�C�sObs��:�ܳ��o��M����X<�8��tLB�B�4���l�2	7� ����17�D,퟉V�m�h���My�O�W��Q��� �b��S"e��_Q�Mj�]dy��f��*���t�M0wV�4pC䓑�R�#���(���+$���$c�
.4����h�v0�9�确i�ε���׊�E�fx�����@���Z��w�+��$���0�	W�P`��Ih��X9��q%	�/$u�$���!��NXnc�����(f��cYy�ˠ�%��lv���Cm�._Q����P��`d����� ʭs��!m�E��{і�a$IY߁ ����@m]UŏV��C���&�Nٱ���p��6����O}F����G��BzG<��W���F�C�>����L�&�m���37Ѳ�=��It.��X:�nA��Gc��/�be`��8%Ĕs��*�(x�����؍"��1r�غ�dĐ � ёO�Ma�R����B[�R^IVZ* ��p��.֡��}�P�F58X����2X�n.Q�o70/�!)�f|��q�e�4� m���������@`�e<���/؛wZ{ (ȏhu�&�I��bfjgڭ�8֚0[Z�C!u0f���Iy(�އ���d�L��v��u�GPgO�$���0k�5n���s��Ym��ŏ�L�V�/�!�֙-I!!P%�r�3;�N�M{=Yl����5'��o1����UӉ?:`7�I۷je�F��*�	Y�!>�uF'�w��O��px�6�iC�B��#VH�u�xS݀VF�`RH(�-�Z��.�p�!�_FN