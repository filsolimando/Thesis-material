BZh91AY&SY a9t 9߁py������?��� @`
���l���|��֜������EU�R��O2jy45L�I��4��dS�� iM=I� 4       �$)��Dh�  �  iI��@    h   DS S�&Ҟ���M@�S@ h4�I	���<�M&P�=M�d  hh�V�e."9D=A� � ����w�B�K=��#1	�Y�>���?u�������n~�(t��1�}s`X�e( y5�-��il[���UUTUUEV�P�@�LnHfBT��^����m��pC&��P$�/\���	��b�)l1T8>	��L�.!āz�Z�_�l�`J�2D��iO[��:��t,��B����*
��c����ߌC�eN)���l�� |
�ķ�'�4�����PL��@�.``�.���P�d5.<ꩧ]2�@�u>�|�!� ����i{I{U�]�67@� ��	�cQ	�v:�!Eg8 �]�b5,v40\�lr�v��O��.L���UT}*5oP$#��� &��I$	��T�C�����hu55(Ԭ�����������\�m㉢b��nӮ�Z�*�'W�u��۷͘B�`B!�j��>1C�:�u�q=f$�,�u�J������il�2)�����Q	�v�ա��O�i���GH�������-u��Z�k~�pnR����t�kUGya�����Q���	�1j��dF�� ��02$���6h�Z������k�1�e���/ ��5��6xh��Ft�(�h��9B��US,W��DC�!�sj��y��C0@��A�C	�
a��@u�o%_S3p�v!2�U�K!�!gf��m\��k[j���z/+&����b�i�G7��Ca�"Q6I%����\� �چ�P�)���[��wg18%t�����Z:��l튙�ֳd��7ZNr��90(������������JS�N�P.�
h��\٪�klMƈD�k\��6�ū�cm[k�
�J�Lam�m]q�+k�ڹ$�\Z��� ډ�������ۄa��GL���[�V�&�Y+$�Vm�@�Ed@�|�ޙ�q��3�M{��*�B�~o|��I!�d�)&z9��=]GV=������a����l�B$S�)���|=���"���݊��\څ�� >�8=9$�5ܷ����!��S_�ߛ�n�@��O�BE
��m�!�a����ٿk���:�Bd��RdG�!j�9�S������ �9^=���%���-�缳Ŵ%Ϣ�黂c����ƅ����C "H"@F+C� �Db&,���``����D��AÜ$-�M-s�������һ���Fy�⻔2����tJ�r�(�����0�C�Ej��@�������wyܤԥ��^�sD�����I �$j�g�w(uD/�'.�!C�m��ƙߨ6>��5�S�yT��6�+��	��xx^�P�@v@ܣ砹M��au)��P�
ߥ�����շ�ũ��ޔ���ju�`K�w� ��wQD �<=���UV��K���`q�[ˢ��6���~�p<�����BKha���}~e��w,.���xaB+���?X��};Ƌ�1m`v>"�æ*͊�H>t���jvxi��O�ZQ�СȖ��j��,�I��h3Ck��k�J�q^
8�3I��b"}El���%ST�H�bȁb/��u��@\�UClā3r�P*���M�
]����p`Z1b�z���$�^i+q��&�N�u�����ۼ@%_��y@%� z^�����3���܁�K��h@�BQCC�Bw6c�����"�w<�n!�'����_q�Q9�H�����^a��,�_Y܉#�А�8	�L�{�sP���A����X �&�Yjc��Cv�M��E������(7t�%���`�F��Y���oQ.!�C]�؇T��*�p�s��9E�HQD@��:���%v�lc��UL��,h� @�92�6�9��3o>1fl�f�s��\��(0H����҆�=QGɈ��*v��rl�B'9�QC�;�nh��M��6H���?N(�z����_����(t�@�S��{�.�p� @�r�